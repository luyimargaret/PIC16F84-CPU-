module sfr(
input clock,
input reset,
input en,
input en_DECODE,
input [5:0]IN_opcode,
input [10:0]IN_operand,
input write_en,
input [7:0]IN_ALU,
output reg en_goto=0,
output reg en_call=0,
output reg en_out=0,
output reg en_short_jump=0,
output reg [9:0]OUT_ALU_PC=0,
output reg mem_wei=1,
output reg [7:0]mem_test=0,
output reg ti
);

reg [7:0]mem[0:255];
always@(posedge clock,posedge reset)
begin
	if(reset==1)
		begin
mem[0]<=8'd0;
mem[1]<=8'd0;
mem[2]<=8'd0;
mem[3]<=8'b0011_1000;
mem[4]<=8'd0;
mem[5]<=8'd0;
mem[6]<=8'd0;
mem[7]<=8'd0;
mem[8]<=8'd0;
mem[9]<=8'd0;
mem[10]<=8'd0;
mem[11]<=8'd0;
mem[12]<=8'd0;
mem[13]<=8'd0;
mem[14]<=8'd0;
mem[15]<=8'd0;
mem[16]<=8'd0;
mem[17]<=8'd0;
mem[18]<=8'd0;
mem[19]<=8'd0;
mem[20]<=8'd0;
mem[21]<=8'd0;
mem[22]<=8'd0;
mem[23]<=8'd0;
mem[24]<=8'd0;
mem[25]<=8'd0;
mem[26]<=8'd0;
mem[27]<=8'd0;
mem[28]<=8'd0;
mem[29]<=8'd0;
mem[30]<=8'd0;
mem[31]<=8'd0;
mem[32]<=8'd0;
mem[33]<=8'd0;
mem[34]<=8'd0;
mem[35]<=8'd0;
mem[36]<=8'd0;
mem[37]<=8'd0;
mem[38]<=8'd0;
mem[39]<=8'd0;
mem[40]<=8'd0;
mem[41]<=8'd0;
mem[42]<=8'd0;
mem[43]<=8'd0;
mem[44]<=8'd0;
mem[45]<=8'd0;
mem[46]<=8'd0;
mem[47]<=8'd0;
mem[48]<=8'd0;
mem[49]<=8'd0;
mem[50]<=8'd0;
mem[51]<=8'd0;
mem[52]<=8'd0;
mem[53]<=8'd0;
mem[54]<=8'd0;
mem[55]<=8'd0;
mem[56]<=8'd0;
mem[57]<=8'd0;
mem[58]<=8'd0;
mem[59]<=8'd0;
mem[60]<=8'd0;
mem[61]<=8'd0;
mem[62]<=8'd0;
mem[63]<=8'd0;
mem[64]<=8'd0;
mem[65]<=8'd0;
mem[66]<=8'd0;
mem[67]<=8'd0;
mem[68]<=8'd0;
mem[69]<=8'd0;
mem[70]<=8'd0;
mem[71]<=8'd0;
mem[72]<=8'd0;
mem[73]<=8'd0;
mem[74]<=8'd0;
mem[75]<=8'd0;
mem[76]<=8'd0;
mem[77]<=8'd0;
mem[78]<=8'd0;
mem[79]<=8'd0;
mem[80]<=8'd0;
mem[81]<=8'd0;
mem[82]<=8'd0;
mem[83]<=8'd0;
mem[84]<=8'd0;
mem[85]<=8'd0;
mem[86]<=8'd0;
mem[87]<=8'd0;
mem[88]<=8'd0;
mem[89]<=8'd0;
mem[90]<=8'd0;
mem[91]<=8'd0;
mem[92]<=8'd0;
mem[93]<=8'd0;
mem[94]<=8'd0;
mem[95]<=8'd0;
mem[96]<=8'd0;
mem[97]<=8'd0;
mem[98]<=8'd0;
mem[99]<=8'd0;
mem[100]<=8'd0;
mem[101]<=8'd0;
mem[102]<=8'd0;
mem[103]<=8'd0;
mem[104]<=8'd0;
mem[105]<=8'd0;
mem[106]<=8'd0;
mem[107]<=8'd0;
mem[108]<=8'd0;
mem[109]<=8'd0;
mem[110]<=8'd0;
mem[111]<=8'd0;
mem[112]<=8'd0;
mem[113]<=8'd0;
mem[114]<=8'd0;
mem[115]<=8'd0;
mem[116]<=8'd0;
mem[117]<=8'd0;
mem[118]<=8'd0;
mem[119]<=8'd0;
mem[120]<=8'd0;
mem[121]<=8'd0;
mem[122]<=8'd0;
mem[123]<=8'd0;
mem[124]<=8'd0;
mem[125]<=8'd0;
mem[126]<=8'd0;
mem[127]<=8'd0;
mem[128]<=8'd0;
mem[129]<=8'd255;
mem[130]<=8'd0;
mem[131]<=8'd0;
mem[132]<=8'd0;
mem[133]<=8'd255;
mem[134]<=8'd255;
mem[135]<=8'd0;
mem[136]<=8'd0;
mem[137]<=8'd0;
mem[138]<=8'd0;
mem[139]<=8'd0;
mem[140]<=8'd0;
mem[141]<=8'd0;
mem[142]<=8'd0;
mem[143]<=8'd255;
mem[144]<=8'd0;
mem[145]<=8'd0;
mem[146]<=8'd0;
mem[147]<=8'd0;
mem[148]<=8'd0;
mem[149]<=8'd0;
mem[150]<=8'd0;
mem[151]<=8'd0;
mem[152]<=8'd0;
mem[153]<=8'd0;
mem[154]<=8'd0;
mem[155]<=8'd0;
mem[156]<=8'd0;
mem[157]<=8'd0;
mem[158]<=8'd0;
mem[159]<=8'd0;
mem[160]<=8'd0;
mem[161]<=8'd0;
mem[162]<=8'd0;
mem[163]<=8'd0;
mem[164]<=8'd0;
mem[165]<=8'd0;
mem[166]<=8'd0;
mem[167]<=8'd0;
mem[168]<=8'd0;
mem[169]<=8'd0;
mem[170]<=8'd0;
mem[171]<=8'd0;
mem[172]<=8'd0;
mem[173]<=8'd0;
mem[174]<=8'd0;
mem[175]<=8'd0;
mem[176]<=8'd0;
mem[177]<=8'd0;
mem[178]<=8'd0;
mem[179]<=8'd0;
mem[180]<=8'd0;
mem[181]<=8'd0;
mem[182]<=8'd0;
mem[183]<=8'd0;
mem[184]<=8'd0;
mem[185]<=8'd0;
mem[186]<=8'd0;
mem[187]<=8'd0;
mem[188]<=8'd0;
mem[189]<=8'd0;
mem[190]<=8'd0;
mem[191]<=8'd0;
mem[192]<=8'd0;
mem[193]<=8'd0;
mem[194]<=8'd0;
mem[195]<=8'd0;
mem[196]<=8'd0;
mem[197]<=8'd0;
mem[198]<=8'd0;
mem[199]<=8'd0;
mem[200]<=8'd0;
mem[201]<=8'd0;
mem[202]<=8'd0;
mem[203]<=8'd0;
mem[204]<=8'd0;
mem[205]<=8'd0;
mem[206]<=8'd0;
mem[207]<=8'd0;
mem[208]<=8'd0;
mem[209]<=8'd0;
mem[210]<=8'd0;
mem[211]<=8'd0;
mem[212]<=8'd0;
mem[213]<=8'd0;
mem[214]<=8'd0;
mem[215]<=8'd0;
mem[216]<=8'd0;
mem[217]<=8'd0;
mem[218]<=8'd0;
mem[219]<=8'd0;
mem[220]<=8'd0;
mem[221]<=8'd0;
mem[222]<=8'd0;
mem[223]<=8'd0;
mem[224]<=8'd0;
mem[225]<=8'd0;
mem[226]<=8'd0;
mem[227]<=8'd0;
mem[228]<=8'd0;
mem[229]<=8'd0;
mem[230]<=8'd0;
mem[231]<=8'd0;
mem[232]<=8'd0;
mem[233]<=8'd0;
mem[234]<=8'd0;
mem[235]<=8'd0;
mem[236]<=8'd0;
mem[237]<=8'd0;
mem[238]<=8'd0;
mem[239]<=8'd0;
mem[240]<=8'd0;
mem[241]<=8'd0;
mem[242]<=8'd0;
mem[243]<=8'd0;
mem[244]<=8'd0;
mem[245]<=8'd0;
mem[246]<=8'd0;
mem[247]<=8'd0;
mem[248]<=8'd0;
mem[249]<=8'd0;
mem[250]<=8'd0;
mem[251]<=8'd0;
mem[252]<=8'd0;
mem[253]<=8'd0;
mem[254]<=8'd0;
mem[255]<=8'd0;

		end
	else
		if((en==1)&&(en_DECODE==1))
		begin
			ti<=1;
			if(mem['h03][5]==1)//选择体1
				begin
				if(IN_opcode==6'd1)//1_CALL
				begin
				en_goto<=0;
				en_call<=1;
				en_out<=0;
				en_short_jump<=0;
				OUT_ALU_PC<=IN_operand[9:0];
				end
			else if(IN_opcode==6'd2)//2_GOTO
				begin
				en_goto<=1;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				OUT_ALU_PC<=IN_operand[9:0];
				end
			else if(IN_opcode==6'd3)//3_BCF
				begin
				mem[IN_operand[6:0]+'d128][IN_operand[9:7]]=0;
				mem_wei=mem[IN_operand[6:0]+'d128][IN_operand[9:7]];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd4)//4_BSF
				begin
				mem[IN_operand[6:0]+'d128][IN_operand[9:7]]=1;
				mem_wei=mem[IN_operand[6:0]+'d128][IN_operand[9:7]];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd5)//5_BTFSC
				begin
				if(mem[IN_operand[6:0]+'d128][IN_operand[9:7]]==0)
					en_short_jump<=1;
				else
					en_short_jump<=0;
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				end
			else if(IN_opcode==6'd6)//6_BTFSS
				begin
				if(mem[IN_operand[6:0]+'d128][IN_operand[9:7]]==1)
					en_short_jump<=1;
				else
					en_short_jump<=0;
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				end
			else if(IN_opcode==6'd8)//8_RETLW
				begin
				en_goto<=0;
				en_call<=0;
				en_out<=1;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd11)//11_SUBWF
				begin
				if(write_en==1)
					begin
					mem[IN_operand[6:0]+'d128]=IN_ALU;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				else
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd12)//12_DECF
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128]-'b1;
				else
					begin
					mem[IN_operand[6:0]+'d128]=mem[IN_operand[6:0]+'d128]-'b1;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd13)//13_IORWF
				begin
				if(write_en==1)
					begin
					mem[IN_operand[6:0]+'d128]=IN_ALU;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				else
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd14)//14_ANDWF
				begin
				if(write_en==1)
					begin
					mem[IN_operand[6:0]+'d128]=IN_ALU;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				else
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end		
			else if(IN_opcode==6'd15)//15_XORWF
				begin
				if(write_en==1)
					begin
					mem[IN_operand[6:0]+'d128]=IN_ALU;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				else
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd16)//16_ADDWF
				begin
				if(write_en==1)
					begin
					mem[IN_operand[6:0]+'d128]=IN_ALU;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				else
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd17)//17_MOVF
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128];
				else
					begin
					mem[IN_operand[6:0]+'d128]=mem[IN_operand[6:0]+'d128];
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd18)//18_COMF
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<=~mem[IN_operand[6:0]+'d128];
				else
					begin
					mem[IN_operand[6:0]+'d128]=~mem[IN_operand[6:0]+'d128];
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd19)//19_INCF
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128]+'b1;
				else
					begin
					mem[IN_operand[6:0]+'d128]=mem[IN_operand[6:0]+'d128]+'b1;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd20)//20_DECFSZ
				begin
				if(mem[IN_operand[6:0]+'d128]-'b1==0)
					en_short_jump<=1;
				else
					en_short_jump<=0;
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128]-'b1;
				else
					begin
					mem[IN_operand[6:0]+'d128]=mem[IN_operand[6:0]+'d128]-'b1;
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				end
			else if(IN_opcode==6'd21)//21_RRF
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<={mem[IN_operand[6:0]+'d128][0],mem[IN_operand[6:0]+'d128][7:1]};
				else
					begin
					mem[IN_operand[6:0]+'d128]={mem[IN_operand[6:0]+'d128][0],mem[IN_operand[6:0]+'d128][7:1]};
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd22)//22_RLF
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<={mem[IN_operand[6:0]+'d128][6:0],mem[IN_operand[6:0]+'d128][7]};
				else
					begin
					mem[IN_operand[6:0]+'d128]={mem[IN_operand[6:0]+'d128][6:0],mem[IN_operand[6:0]+'d128][7]};
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd23)//23_SWAP
				begin
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<={mem[IN_operand[6:0]+'d128][3:0],mem[IN_operand[6:0]+'d128][7:4]};
				else
					begin
					mem[IN_operand[6:0]+'d128]={mem[IN_operand[6:0]+'d128][3:0],mem[IN_operand[6:0]+'d128][7:4]};
					mem_test=mem[IN_operand[6:0]+'d128];
					end
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd24)//24_INCFSZ
				begin
				if(mem[IN_operand[6:0]+'d128]+'b1==9'b10000_0000)
					en_short_jump<=1;
				else
					en_short_jump<=0;
				if(IN_operand[7]==0)
					OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]+'d128]+'b1;
				else
					begin
					mem[IN_operand[6:0]+'d128]=mem[IN_operand[6:0]+'d128]+'b1;
					mem_test=mem[IN_operand[6:0]+'d128];
					end	
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				end
			else if(IN_opcode==6'd28)//28_CLRF
				begin
				mem[IN_operand[6:0]+'d128]=0;
				mem_test=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd30)//30_MOVWF
				begin
				mem[IN_operand[6:0]+'d128]=IN_ALU;
				mem_test=mem[IN_operand[6:0]+'d128];
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd32)//32_RETURN	
				begin
				en_goto<=0;
				en_call<=0;
				en_out<=1;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd33)//33_RETFIE	
				begin
				mem['h0b+'d128][7]=1'b1;
				mem_wei=mem['h0b+'d128][7];
				en_goto<=0;
				en_call<=0;
				en_out<=1;
				en_short_jump<=0;
				end
			else if(IN_opcode==6'd34)//34_SLEEP	
				begin
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else if(IN_opcode==6'd35)//35_CLRWDT
				begin
				en_goto<=0;
				en_call<=0;
				en_out<=0;
				en_short_jump<=0;
				end	
			else
				begin
				en_goto<=en_goto;
				en_call<=en_call;
				en_out<=en_out;
				en_short_jump<=en_short_jump;
				OUT_ALU_PC<=OUT_ALU_PC;
				mem_wei<=mem_wei;
				mem_test<=mem_test;
				end
				end
///////////////////////////////////////////////////////////////////////				
			else//选择体0
				begin
				ti<=0;
				if(IN_opcode==6'd1)//1_CALL
					begin
					en_goto<=0;
					en_call<=1;
					en_out<=0;
					en_short_jump<=0;
					OUT_ALU_PC<=IN_operand[9:0];
					end
				else if(IN_opcode==6'd2)//2_GOTO
					begin
					en_goto<=1;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					OUT_ALU_PC<=IN_operand[9:0];
					end
				else if(IN_opcode==6'd3)//3_BCF
					begin
					mem[IN_operand[6:0]][IN_operand[9:7]]=0;
					mem_wei=mem[IN_operand[6:0]][IN_operand[9:7]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd4)//4_BSF
					begin	
					mem[IN_operand[6:0]][IN_operand[9:7]]=1;
					mem_wei=mem[IN_operand[6:0]][IN_operand[9:7]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd5)//5_BTFSC
					begin
					if(mem[IN_operand[6:0]][IN_operand[9:7]]==0)
						en_short_jump<=1;
					else
						en_short_jump<=0;
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					end
				else if(IN_opcode==6'd6)//6_BTFSS
					begin
					if(mem[IN_operand[6:0]][IN_operand[9:7]]==1)
						en_short_jump<=1;
					else
						en_short_jump<=0;
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					end
				else if(IN_opcode==6'd8)//8_RETLW
					begin
					en_goto<=0;
					en_call<=0;
					en_out<=1;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd11)//11_SUBWF
					begin
					if(write_en==1)
						begin
						mem[IN_operand[6:0]]=IN_ALU;
						mem_test=mem[IN_operand[6:0]];
						end
					else
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd12)//12_DECF
					begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]]-'b1;
					else
						begin
						mem[IN_operand[6:0]]=mem[IN_operand[6:0]]-'b1;
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd13)//13_IORWF
					begin
					if(write_en==1)
					begin
						mem[IN_operand[6:0]]=IN_ALU;
						mem_test=mem[IN_operand[6:0]];
						end
					else
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd14)//14_ANDWF
					begin
					if(write_en==1)
					begin
						mem[IN_operand[6:0]]=IN_ALU;
						mem_test=mem[IN_operand[6:0]];
					end
					else
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end		
				else if(IN_opcode==6'd15)//15_XORWF
					begin
					if(write_en==1)
						begin
						mem[IN_operand[6:0]]=IN_ALU;
						mem_test=mem[IN_operand[6:0]];
						end
					else
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd16)//16_ADDWF
					begin
					if(write_en==1)
						begin
						mem[IN_operand[6:0]]=IN_ALU;
						mem_test=mem[IN_operand[6:0]];
						end
					else
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd17)//17_MOVF
					begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]];
					else
						begin
						mem[IN_operand[6:0]]=mem[IN_operand[6:0]];
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd18)//18_COMF
					begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<=~mem[IN_operand[6:0]];
					else
						begin
						mem[IN_operand[6:0]]=~mem[IN_operand[6:0]];
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd19)//19_INCF
					begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]]+'b1;
					else
						begin
						mem[IN_operand[6:0]]=mem[IN_operand[6:0]]+'b1;
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd20)//20_DECFSZ
					begin
					if(mem[IN_operand[6:0]]-'b1==0)
						en_short_jump<=1;
					else
						en_short_jump<=0;
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]]-'b1;
					else
						begin
						mem[IN_operand[6:0]]=mem[IN_operand[6:0]]-'b1;
						mem_test=mem[IN_operand[6:0]];
						end	
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					end
				else if(IN_opcode==6'd21)//21_RRF
					begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<={mem[IN_operand[6:0]][0],mem[IN_operand[6:0]][7:1]};
					else
						begin
						mem[IN_operand[6:0]]={mem[IN_operand[6:0]][0],mem[IN_operand[6:0]][7:1]};
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd22)//22_RLF
				begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<={mem[IN_operand[6:0]][6:0],mem[IN_operand[6:0]][7]};
					else
						begin
						mem[IN_operand[6:0]]={mem[IN_operand[6:0]][6:0],mem[IN_operand[6:0]][7]};
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd23)//23_SWAP
					begin
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<={mem[IN_operand[6:0]][3:0],mem[IN_operand[6:0]][7:4]};
					else
						begin
						mem[IN_operand[6:0]]={mem[IN_operand[6:0]][3:0],mem[IN_operand[6:0]][7:4]};
						mem_test=mem[IN_operand[6:0]];
						end
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd24)//24_INCFSZ
					begin
					if(mem[IN_operand[6:0]]+'b1==9'b10000_0000)
						en_short_jump<=1;
					else
						en_short_jump<=0;
					if(IN_operand[7]==0)
						OUT_ALU_PC[7:0]<=mem[IN_operand[6:0]]+'b1;
					else
						begin
						mem[IN_operand[6:0]]=mem[IN_operand[6:0]]+'b1;
						mem_test=mem[IN_operand[6:0]];
						end	
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					end
				else if(IN_opcode==6'd28)//28_CLRF
					begin
						mem[IN_operand[6:0]]=0;
						mem_test=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd30)//30_MOVWF
					begin
					mem[IN_operand[6:0]]=IN_ALU;
					mem_test=mem[IN_operand[6:0]];
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd32)//32_RETURN	
					begin
					en_goto<=0;
					en_call<=0;
					en_out<=1;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd33)//33_RETFIE	
					begin
					mem['h0b][7]=1'b1;
					mem_wei=mem['h0b][7];
					en_goto<=0;
					en_call<=0;
					en_out<=1;
					en_short_jump<=0;
					end
				else if(IN_opcode==6'd34)//34_SLEEP	
					begin
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else if(IN_opcode==6'd35)//35_CLRWDT
					begin
					en_goto<=0;
					en_call<=0;
					en_out<=0;
					en_short_jump<=0;
					end	
				else
					begin
					en_goto<=en_goto;
					en_call<=en_call;
					en_out<=en_out;
					en_short_jump<=en_short_jump;
					OUT_ALU_PC<=OUT_ALU_PC;
					mem_wei<=mem_wei;
					mem_test<=mem_test;
					end
				end//end选择体0的else
			end//end的是if(en&&en_DECODE)
		else
			begin
			en_goto<=en_goto;
			en_call<=en_call;
			en_out<=en_out;
			en_short_jump<=en_short_jump;
			OUT_ALU_PC<=OUT_ALU_PC;
			mem_wei<=mem_wei;
			mem_test<=mem_test;
			end
end//end的是always开始的begin
endmodule


