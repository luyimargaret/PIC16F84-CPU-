module memory(
input clock,
input reset,
input[9:0]IN_PC,
input en,
output reg[13:0]OUT_DECODE=0
);

reg[13:0]mem[0:1023];

always@(posedge clock,posedge reset)
begin
	if(reset==1)
		begin
mem[0]<='h0183;
mem[1]<='h3000;
mem[2]<='h008A;
mem[3]<='h2804;
mem[4]<='h0183;
mem[5]<='h3003;
mem[6]<='h00AD;
mem[7]<='h30E7;
mem[8]<='h00AC;
mem[9]<='h3012;
mem[10]<='h0084;
mem[11]<='h302B;
mem[12]<='h200F;
mem[13]<='h0183;
mem[14]<='h2B91;
mem[15]<='h00AB;
mem[16]<='h201A;
mem[17]<='h0080;
mem[18]<='h0A84;
mem[19]<='h0804;
mem[20]<='h062B;
mem[21]<='h1903;
mem[22]<='h3400;
mem[23]<='h2810;
mem[24]<='h1283;
mem[25]<='h00AC;
mem[26]<='h1BAD;
mem[27]<='h2823;
mem[28]<='h082D;
mem[29]<='h008A;
mem[30]<='h082C;
mem[31]<='h0AAC;
mem[32]<='h1903;
mem[33]<='h0AAD;
mem[34]<='h0082;
mem[35]<='h1383;
mem[36]<='h182D;
mem[37]<='h1783;
mem[38]<='h082C;
mem[39]<='h0AAC;
mem[40]<='h0084;
mem[41]<='h0800;
mem[42]<='h0008;
mem[43]<='h3fff;
mem[44]<='h3fff;
mem[45]<='h3fff;
mem[46]<='h3fff;
mem[47]<='h3fff;
mem[48]<='h3fff;
mem[49]<='h3fff;
mem[50]<='h3fff;
mem[51]<='h3fff;
mem[52]<='h3fff;
mem[53]<='h3fff;
mem[54]<='h3fff;
mem[55]<='h3fff;
mem[56]<='h3fff;
mem[57]<='h3fff;
mem[58]<='h3fff;
mem[59]<='h3fff;
mem[60]<='h3fff;
mem[61]<='h3fff;
mem[62]<='h3fff;
mem[63]<='h3fff;
mem[64]<='h3fff;
mem[65]<='h3fff;
mem[66]<='h3fff;
mem[67]<='h3fff;
mem[68]<='h3fff;
mem[69]<='h3fff;
mem[70]<='h3fff;
mem[71]<='h3fff;
mem[72]<='h3fff;
mem[73]<='h3fff;
mem[74]<='h3fff;
mem[75]<='h3fff;
mem[76]<='h3fff;
mem[77]<='h3fff;
mem[78]<='h3fff;
mem[79]<='h3fff;
mem[80]<='h3fff;
mem[81]<='h3fff;
mem[82]<='h3fff;
mem[83]<='h3fff;
mem[84]<='h3fff;
mem[85]<='h3fff;
mem[86]<='h3fff;
mem[87]<='h3fff;
mem[88]<='h3fff;
mem[89]<='h3fff;
mem[90]<='h3fff;
mem[91]<='h3fff;
mem[92]<='h3fff;
mem[93]<='h3fff;
mem[94]<='h3fff;
mem[95]<='h3fff;
mem[96]<='h3fff;
mem[97]<='h3fff;
mem[98]<='h3fff;
mem[99]<='h3fff;
mem[100]<='h3fff;
mem[101]<='h3fff;
mem[102]<='h3fff;
mem[103]<='h3fff;
mem[104]<='h3fff;
mem[105]<='h3fff;
mem[106]<='h3fff;
mem[107]<='h3fff;
mem[108]<='h3fff;
mem[109]<='h3fff;
mem[110]<='h3fff;
mem[111]<='h3fff;
mem[112]<='h3fff;
mem[113]<='h3fff;
mem[114]<='h3fff;
mem[115]<='h3fff;
mem[116]<='h3fff;
mem[117]<='h3fff;
mem[118]<='h3fff;
mem[119]<='h3fff;
mem[120]<='h3fff;
mem[121]<='h3fff;
mem[122]<='h3fff;
mem[123]<='h3fff;
mem[124]<='h3fff;
mem[125]<='h3fff;
mem[126]<='h3fff;
mem[127]<='h3fff;
mem[128]<='h3fff;
mem[129]<='h3fff;
mem[130]<='h3fff;
mem[131]<='h3fff;
mem[132]<='h3fff;
mem[133]<='h3fff;
mem[134]<='h3fff;
mem[135]<='h3fff;
mem[136]<='h3fff;
mem[137]<='h3fff;
mem[138]<='h3fff;
mem[139]<='h3fff;
mem[140]<='h3fff;
mem[141]<='h3fff;
mem[142]<='h3fff;
mem[143]<='h3fff;
mem[144]<='h3fff;
mem[145]<='h3fff;
mem[146]<='h3fff;
mem[147]<='h3fff;
mem[148]<='h3fff;
mem[149]<='h3fff;
mem[150]<='h3fff;
mem[151]<='h3fff;
mem[152]<='h3fff;
mem[153]<='h3fff;
mem[154]<='h3fff;
mem[155]<='h3fff;
mem[156]<='h3fff;
mem[157]<='h3fff;
mem[158]<='h3fff;
mem[159]<='h3fff;
mem[160]<='h3fff;
mem[161]<='h3fff;
mem[162]<='h3fff;
mem[163]<='h3fff;
mem[164]<='h3fff;
mem[165]<='h3fff;
mem[166]<='h3fff;
mem[167]<='h3fff;
mem[168]<='h3fff;
mem[169]<='h3fff;
mem[170]<='h3fff;
mem[171]<='h3fff;
mem[172]<='h3fff;
mem[173]<='h3fff;
mem[174]<='h3fff;
mem[175]<='h3fff;
mem[176]<='h3fff;
mem[177]<='h3fff;
mem[178]<='h3fff;
mem[179]<='h3fff;
mem[180]<='h3fff;
mem[181]<='h3fff;
mem[182]<='h3fff;
mem[183]<='h3fff;
mem[184]<='h3fff;
mem[185]<='h3fff;
mem[186]<='h3fff;
mem[187]<='h3fff;
mem[188]<='h3fff;
mem[189]<='h3fff;
mem[190]<='h3fff;
mem[191]<='h3fff;
mem[192]<='h3fff;
mem[193]<='h3fff;
mem[194]<='h3fff;
mem[195]<='h3fff;
mem[196]<='h3fff;
mem[197]<='h3fff;
mem[198]<='h3fff;
mem[199]<='h3fff;
mem[200]<='h3fff;
mem[201]<='h3fff;
mem[202]<='h3fff;
mem[203]<='h3fff;
mem[204]<='h3fff;
mem[205]<='h3fff;
mem[206]<='h3fff;
mem[207]<='h3fff;
mem[208]<='h3fff;
mem[209]<='h3fff;
mem[210]<='h3fff;
mem[211]<='h3fff;
mem[212]<='h3fff;
mem[213]<='h3fff;
mem[214]<='h3fff;
mem[215]<='h3fff;
mem[216]<='h3fff;
mem[217]<='h3fff;
mem[218]<='h3fff;
mem[219]<='h3fff;
mem[220]<='h3fff;
mem[221]<='h3fff;
mem[222]<='h3fff;
mem[223]<='h3fff;
mem[224]<='h3fff;
mem[225]<='h3fff;
mem[226]<='h3fff;
mem[227]<='h3fff;
mem[228]<='h3fff;
mem[229]<='h3fff;
mem[230]<='h3fff;
mem[231]<='h3fff;
mem[232]<='h3fff;
mem[233]<='h3fff;
mem[234]<='h3fff;
mem[235]<='h3fff;
mem[236]<='h3fff;
mem[237]<='h3fff;
mem[238]<='h3fff;
mem[239]<='h3fff;
mem[240]<='h3fff;
mem[241]<='h3fff;
mem[242]<='h3fff;
mem[243]<='h3fff;
mem[244]<='h3fff;
mem[245]<='h3fff;
mem[246]<='h3fff;
mem[247]<='h3fff;
mem[248]<='h3fff;
mem[249]<='h3fff;
mem[250]<='h3fff;
mem[251]<='h3fff;
mem[252]<='h3fff;
mem[253]<='h3fff;
mem[254]<='h3fff;
mem[255]<='h3fff;
mem[256]<='h3fff;
mem[257]<='h3fff;
mem[258]<='h3fff;
mem[259]<='h3fff;
mem[260]<='h3fff;
mem[261]<='h3fff;
mem[262]<='h3fff;
mem[263]<='h3fff;
mem[264]<='h3fff;
mem[265]<='h3fff;
mem[266]<='h3fff;
mem[267]<='h3fff;
mem[268]<='h3fff;
mem[269]<='h3fff;
mem[270]<='h3fff;
mem[271]<='h3fff;
mem[272]<='h3fff;
mem[273]<='h3fff;
mem[274]<='h3fff;
mem[275]<='h3fff;
mem[276]<='h3fff;
mem[277]<='h3fff;
mem[278]<='h3fff;
mem[279]<='h3fff;
mem[280]<='h3fff;
mem[281]<='h3fff;
mem[282]<='h3fff;
mem[283]<='h3fff;
mem[284]<='h3fff;
mem[285]<='h3fff;
mem[286]<='h3fff;
mem[287]<='h3fff;
mem[288]<='h3fff;
mem[289]<='h3fff;
mem[290]<='h3fff;
mem[291]<='h3fff;
mem[292]<='h3fff;
mem[293]<='h3fff;
mem[294]<='h3fff;
mem[295]<='h3fff;
mem[296]<='h3fff;
mem[297]<='h3fff;
mem[298]<='h3fff;
mem[299]<='h3fff;
mem[300]<='h3fff;
mem[301]<='h3fff;
mem[302]<='h3fff;
mem[303]<='h3fff;
mem[304]<='h3fff;
mem[305]<='h3fff;
mem[306]<='h3fff;
mem[307]<='h3fff;
mem[308]<='h3fff;
mem[309]<='h3fff;
mem[310]<='h3fff;
mem[311]<='h3fff;
mem[312]<='h3fff;
mem[313]<='h3fff;
mem[314]<='h3fff;
mem[315]<='h3fff;
mem[316]<='h3fff;
mem[317]<='h3fff;
mem[318]<='h3fff;
mem[319]<='h3fff;
mem[320]<='h3fff;
mem[321]<='h3fff;
mem[322]<='h3fff;
mem[323]<='h3fff;
mem[324]<='h3fff;
mem[325]<='h3fff;
mem[326]<='h3fff;
mem[327]<='h3fff;
mem[328]<='h3fff;
mem[329]<='h3fff;
mem[330]<='h3fff;
mem[331]<='h3fff;
mem[332]<='h3fff;
mem[333]<='h3fff;
mem[334]<='h3fff;
mem[335]<='h3fff;
mem[336]<='h3fff;
mem[337]<='h3fff;
mem[338]<='h3fff;
mem[339]<='h3fff;
mem[340]<='h3fff;
mem[341]<='h3fff;
mem[342]<='h3fff;
mem[343]<='h3fff;
mem[344]<='h3fff;
mem[345]<='h3fff;
mem[346]<='h3fff;
mem[347]<='h3fff;
mem[348]<='h3fff;
mem[349]<='h3fff;
mem[350]<='h3fff;
mem[351]<='h3fff;
mem[352]<='h3fff;
mem[353]<='h3fff;
mem[354]<='h3fff;
mem[355]<='h3fff;
mem[356]<='h3fff;
mem[357]<='h3fff;
mem[358]<='h3fff;
mem[359]<='h3fff;
mem[360]<='h3fff;
mem[361]<='h3fff;
mem[362]<='h3fff;
mem[363]<='h3fff;
mem[364]<='h3fff;
mem[365]<='h3fff;
mem[366]<='h3fff;
mem[367]<='h3fff;
mem[368]<='h3fff;
mem[369]<='h3fff;
mem[370]<='h3fff;
mem[371]<='h3fff;
mem[372]<='h3fff;
mem[373]<='h3fff;
mem[374]<='h3fff;
mem[375]<='h3fff;
mem[376]<='h3fff;
mem[377]<='h3fff;
mem[378]<='h3fff;
mem[379]<='h3fff;
mem[380]<='h3fff;
mem[381]<='h3fff;
mem[382]<='h3fff;
mem[383]<='h3fff;
mem[384]<='h3fff;
mem[385]<='h3fff;
mem[386]<='h3fff;
mem[387]<='h3fff;
mem[388]<='h3fff;
mem[389]<='h3fff;
mem[390]<='h3fff;
mem[391]<='h3fff;
mem[392]<='h3fff;
mem[393]<='h3fff;
mem[394]<='h3fff;
mem[395]<='h3fff;
mem[396]<='h3fff;
mem[397]<='h3fff;
mem[398]<='h3fff;
mem[399]<='h3fff;
mem[400]<='h3fff;
mem[401]<='h3fff;
mem[402]<='h3fff;
mem[403]<='h3fff;
mem[404]<='h3fff;
mem[405]<='h3fff;
mem[406]<='h3fff;
mem[407]<='h3fff;
mem[408]<='h3fff;
mem[409]<='h3fff;
mem[410]<='h3fff;
mem[411]<='h3fff;
mem[412]<='h3fff;
mem[413]<='h3fff;
mem[414]<='h3fff;
mem[415]<='h3fff;
mem[416]<='h3fff;
mem[417]<='h3fff;
mem[418]<='h3fff;
mem[419]<='h3fff;
mem[420]<='h3fff;
mem[421]<='h3fff;
mem[422]<='h3fff;
mem[423]<='h3fff;
mem[424]<='h3fff;
mem[425]<='h3fff;
mem[426]<='h3fff;
mem[427]<='h3fff;
mem[428]<='h3fff;
mem[429]<='h3fff;
mem[430]<='h3fff;
mem[431]<='h3fff;
mem[432]<='h3fff;
mem[433]<='h3fff;
mem[434]<='h3fff;
mem[435]<='h3fff;
mem[436]<='h3fff;
mem[437]<='h3fff;
mem[438]<='h3fff;
mem[439]<='h3fff;
mem[440]<='h3fff;
mem[441]<='h3fff;
mem[442]<='h3fff;
mem[443]<='h3fff;
mem[444]<='h3fff;
mem[445]<='h3fff;
mem[446]<='h3fff;
mem[447]<='h3fff;
mem[448]<='h3fff;
mem[449]<='h3fff;
mem[450]<='h3fff;
mem[451]<='h3fff;
mem[452]<='h3fff;
mem[453]<='h3fff;
mem[454]<='h3fff;
mem[455]<='h3fff;
mem[456]<='h3fff;
mem[457]<='h3fff;
mem[458]<='h3fff;
mem[459]<='h3fff;
mem[460]<='h3fff;
mem[461]<='h3fff;
mem[462]<='h3fff;
mem[463]<='h3fff;
mem[464]<='h3fff;
mem[465]<='h3fff;
mem[466]<='h3fff;
mem[467]<='h3fff;
mem[468]<='h3fff;
mem[469]<='h3fff;
mem[470]<='h3fff;
mem[471]<='h3fff;
mem[472]<='h3fff;
mem[473]<='h3fff;
mem[474]<='h3fff;
mem[475]<='h3fff;
mem[476]<='h3fff;
mem[477]<='h3fff;
mem[478]<='h3fff;
mem[479]<='h3fff;
mem[480]<='h3fff;
mem[481]<='h3fff;
mem[482]<='h3fff;
mem[483]<='h3fff;
mem[484]<='h3fff;
mem[485]<='h3fff;
mem[486]<='h3fff;
mem[487]<='h3fff;
mem[488]<='h3fff;
mem[489]<='h3fff;
mem[490]<='h3fff;
mem[491]<='h3fff;
mem[492]<='h3fff;
mem[493]<='h3fff;
mem[494]<='h3fff;
mem[495]<='h3fff;
mem[496]<='h3fff;
mem[497]<='h3fff;
mem[498]<='h3fff;
mem[499]<='h3fff;
mem[500]<='h3fff;
mem[501]<='h3fff;
mem[502]<='h3fff;
mem[503]<='h3fff;
mem[504]<='h3fff;
mem[505]<='h3fff;
mem[506]<='h3fff;
mem[507]<='h3fff;
mem[508]<='h3fff;
mem[509]<='h3fff;
mem[510]<='h3fff;
mem[511]<='h3fff;
mem[512]<='h3fff;
mem[513]<='h3fff;
mem[514]<='h3fff;
mem[515]<='h3fff;
mem[516]<='h3fff;
mem[517]<='h3fff;
mem[518]<='h3fff;
mem[519]<='h3fff;
mem[520]<='h3fff;
mem[521]<='h3fff;
mem[522]<='h3fff;
mem[523]<='h3fff;
mem[524]<='h3fff;
mem[525]<='h3fff;
mem[526]<='h3fff;
mem[527]<='h3fff;
mem[528]<='h3fff;
mem[529]<='h3fff;
mem[530]<='h3fff;
mem[531]<='h3fff;
mem[532]<='h3fff;
mem[533]<='h3fff;
mem[534]<='h3fff;
mem[535]<='h3fff;
mem[536]<='h3fff;
mem[537]<='h3fff;
mem[538]<='h3fff;
mem[539]<='h3fff;
mem[540]<='h3fff;
mem[541]<='h3fff;
mem[542]<='h3fff;
mem[543]<='h3fff;
mem[544]<='h3fff;
mem[545]<='h3fff;
mem[546]<='h3fff;
mem[547]<='h3fff;
mem[548]<='h3fff;
mem[549]<='h3fff;
mem[550]<='h3fff;
mem[551]<='h3fff;
mem[552]<='h3fff;
mem[553]<='h3fff;
mem[554]<='h3fff;
mem[555]<='h3fff;
mem[556]<='h3fff;
mem[557]<='h3fff;
mem[558]<='h3fff;
mem[559]<='h3fff;
mem[560]<='h3fff;
mem[561]<='h3fff;
mem[562]<='h3fff;
mem[563]<='h3fff;
mem[564]<='h3fff;
mem[565]<='h3fff;
mem[566]<='h3fff;
mem[567]<='h3fff;
mem[568]<='h3fff;
mem[569]<='h3fff;
mem[570]<='h3fff;
mem[571]<='h3fff;
mem[572]<='h3fff;
mem[573]<='h3fff;
mem[574]<='h3fff;
mem[575]<='h3fff;
mem[576]<='h3fff;
mem[577]<='h3fff;
mem[578]<='h3fff;
mem[579]<='h3fff;
mem[580]<='h3fff;
mem[581]<='h3fff;
mem[582]<='h3fff;
mem[583]<='h3fff;
mem[584]<='h3fff;
mem[585]<='h3fff;
mem[586]<='h3fff;
mem[587]<='h3fff;
mem[588]<='h3fff;
mem[589]<='h3fff;
mem[590]<='h3fff;
mem[591]<='h3fff;
mem[592]<='h3fff;
mem[593]<='h3fff;
mem[594]<='h3fff;
mem[595]<='h3fff;
mem[596]<='h3fff;
mem[597]<='h3fff;
mem[598]<='h3fff;
mem[599]<='h3fff;
mem[600]<='h3fff;
mem[601]<='h3fff;
mem[602]<='h3fff;
mem[603]<='h3fff;
mem[604]<='h3fff;
mem[605]<='h3fff;
mem[606]<='h3fff;
mem[607]<='h3fff;
mem[608]<='h3fff;
mem[609]<='h3fff;
mem[610]<='h3fff;
mem[611]<='h3fff;
mem[612]<='h3fff;
mem[613]<='h3fff;
mem[614]<='h3fff;
mem[615]<='h3fff;
mem[616]<='h3fff;
mem[617]<='h3fff;
mem[618]<='h3fff;
mem[619]<='h3fff;
mem[620]<='h3fff;
mem[621]<='h3fff;
mem[622]<='h3fff;
mem[623]<='h3fff;
mem[624]<='h3fff;
mem[625]<='h3fff;
mem[626]<='h3fff;
mem[627]<='h3fff;
mem[628]<='h3fff;
mem[629]<='h3fff;
mem[630]<='h3fff;
mem[631]<='h3fff;
mem[632]<='h3fff;
mem[633]<='h3fff;
mem[634]<='h3fff;
mem[635]<='h3fff;
mem[636]<='h3fff;
mem[637]<='h3fff;
mem[638]<='h3fff;
mem[639]<='h3fff;
mem[640]<='h3fff;
mem[641]<='h3fff;
mem[642]<='h3fff;
mem[643]<='h3fff;
mem[644]<='h3fff;
mem[645]<='h3fff;
mem[646]<='h3fff;
mem[647]<='h3fff;
mem[648]<='h3fff;
mem[649]<='h3fff;
mem[650]<='h3fff;
mem[651]<='h3fff;
mem[652]<='h3fff;
mem[653]<='h3fff;
mem[654]<='h3fff;
mem[655]<='h3fff;
mem[656]<='h3fff;
mem[657]<='h3fff;
mem[658]<='h3fff;
mem[659]<='h3fff;
mem[660]<='h3fff;
mem[661]<='h3fff;
mem[662]<='h3fff;
mem[663]<='h3fff;
mem[664]<='h3fff;
mem[665]<='h3fff;
mem[666]<='h3fff;
mem[667]<='h3fff;
mem[668]<='h3fff;
mem[669]<='h3fff;
mem[670]<='h3fff;
mem[671]<='h3fff;
mem[672]<='h3fff;
mem[673]<='h3fff;
mem[674]<='h3fff;
mem[675]<='h3fff;
mem[676]<='h3fff;
mem[677]<='h3fff;
mem[678]<='h3fff;
mem[679]<='h3fff;
mem[680]<='h3fff;
mem[681]<='h3fff;
mem[682]<='h3fff;
mem[683]<='h3fff;
mem[684]<='h3fff;
mem[685]<='h3fff;
mem[686]<='h3fff;
mem[687]<='h3fff;
mem[688]<='h3fff;
mem[689]<='h3fff;
mem[690]<='h3fff;
mem[691]<='h3fff;
mem[692]<='h3fff;
mem[693]<='h3fff;
mem[694]<='h3fff;
mem[695]<='h3fff;
mem[696]<='h3fff;
mem[697]<='h3fff;
mem[698]<='h3fff;
mem[699]<='h3fff;
mem[700]<='h3fff;
mem[701]<='h3fff;
mem[702]<='h3fff;
mem[703]<='h3fff;
mem[704]<='h3fff;
mem[705]<='h3fff;
mem[706]<='h3fff;
mem[707]<='h3fff;
mem[708]<='h3fff;
mem[709]<='h3fff;
mem[710]<='h3fff;
mem[711]<='h3fff;
mem[712]<='h3fff;
mem[713]<='h3fff;
mem[714]<='h3fff;
mem[715]<='h3fff;
mem[716]<='h3fff;
mem[717]<='h3fff;
mem[718]<='h3fff;
mem[719]<='h3fff;
mem[720]<='h3fff;
mem[721]<='h3fff;
mem[722]<='h3fff;
mem[723]<='h3fff;
mem[724]<='h3fff;
mem[725]<='h3fff;
mem[726]<='h3fff;
mem[727]<='h3fff;
mem[728]<='h3fff;
mem[729]<='h3fff;
mem[730]<='h3fff;
mem[731]<='h3fff;
mem[732]<='h3fff;
mem[733]<='h3fff;
mem[734]<='h3fff;
mem[735]<='h3fff;
mem[736]<='h3fff;
mem[737]<='h3fff;
mem[738]<='h3fff;
mem[739]<='h3fff;
mem[740]<='h3fff;
mem[741]<='h3fff;
mem[742]<='h3fff;
mem[743]<='h3fff;
mem[744]<='h3fff;
mem[745]<='h3fff;
mem[746]<='h3fff;
mem[747]<='h3fff;
mem[748]<='h3fff;
mem[749]<='h3fff;
mem[750]<='h3fff;
mem[751]<='h3fff;
mem[752]<='h3fff;
mem[753]<='h3fff;
mem[754]<='h3fff;
mem[755]<='h3fff;
mem[756]<='h3fff;
mem[757]<='h3fff;
mem[758]<='h3fff;
mem[759]<='h3fff;
mem[760]<='h3fff;
mem[761]<='h3fff;
mem[762]<='h3fff;
mem[763]<='h3fff;
mem[764]<='h3fff;
mem[765]<='h3fff;
mem[766]<='h3fff;
mem[767]<='h3fff;
mem[768]<='h3fff;
mem[769]<='h3fff;
mem[770]<='h3fff;
mem[771]<='h3fff;
mem[772]<='h3fff;
mem[773]<='h3fff;
mem[774]<='h3fff;
mem[775]<='h3fff;
mem[776]<='h3fff;
mem[777]<='h3fff;
mem[778]<='h3fff;
mem[779]<='h3fff;
mem[780]<='h3fff;
mem[781]<='h3fff;
mem[782]<='h3fff;
mem[783]<='h3fff;
mem[784]<='h3fff;
mem[785]<='h3fff;
mem[786]<='h3fff;
mem[787]<='h3fff;
mem[788]<='h3fff;
mem[789]<='h3fff;
mem[790]<='h3fff;
mem[791]<='h3fff;
mem[792]<='h3fff;
mem[793]<='h3fff;
mem[794]<='h3fff;
mem[795]<='h3fff;
mem[796]<='h3fff;
mem[797]<='h3fff;
mem[798]<='h3fff;
mem[799]<='h3fff;
mem[800]<='h3fff;
mem[801]<='h3fff;
mem[802]<='h3fff;
mem[803]<='h3fff;
mem[804]<='h3fff;
mem[805]<='h3fff;
mem[806]<='h3fff;
mem[807]<='h3fff;
mem[808]<='h3fff;
mem[809]<='h3fff;
mem[810]<='h3fff;
mem[811]<='h3fff;
mem[812]<='h3fff;
mem[813]<='h3fff;
mem[814]<='h3fff;
mem[815]<='h3fff;
mem[816]<='h3fff;
mem[817]<='h3fff;
mem[818]<='h3fff;
mem[819]<='h3fff;
mem[820]<='h3fff;
mem[821]<='h3fff;
mem[822]<='h3fff;
mem[823]<='h3fff;
mem[824]<='h3fff;
mem[825]<='h3fff;
mem[826]<='h3fff;
mem[827]<='h3fff;
mem[828]<='h3fff;
mem[829]<='h3fff;
mem[830]<='h3fff;
mem[831]<='h3fff;
mem[832]<='h3fff;
mem[833]<='h3fff;
mem[834]<='h3fff;
mem[835]<='h3fff;
mem[836]<='h3fff;
mem[837]<='h3fff;
mem[838]<='h3fff;
mem[839]<='h3fff;
mem[840]<='h3fff;
mem[841]<='h3fff;
mem[842]<='h3fff;
mem[843]<='h3fff;
mem[844]<='h3fff;
mem[845]<='h3fff;
mem[846]<='h3fff;
mem[847]<='h3fff;
mem[848]<='h3fff;
mem[849]<='h3fff;
mem[850]<='h3fff;
mem[851]<='h3fff;
mem[852]<='h3fff;
mem[853]<='h3fff;
mem[854]<='h3fff;
mem[855]<='h3fff;
mem[856]<='h3fff;
mem[857]<='h3fff;
mem[858]<='h3fff;
mem[859]<='h3fff;
mem[860]<='h3fff;
mem[861]<='h3fff;
mem[862]<='h3fff;
mem[863]<='h3fff;
mem[864]<='h3fff;
mem[865]<='h3fff;
mem[866]<='h3fff;
mem[867]<='h3fff;
mem[868]<='h3fff;
mem[869]<='h3fff;
mem[870]<='h3fff;
mem[871]<='h3fff;
mem[872]<='h3fff;
mem[873]<='h3fff;
mem[874]<='h3fff;
mem[875]<='h3fff;
mem[876]<='h3fff;
mem[877]<='h3fff;
mem[878]<='h3fff;
mem[879]<='h3fff;
mem[880]<='h3fff;
mem[881]<='h3fff;
mem[882]<='h3fff;
mem[883]<='h3fff;
mem[884]<='h3fff;
mem[885]<='h3fff;
mem[886]<='h3fff;
mem[887]<='h3fff;
mem[888]<='h3fff;
mem[889]<='h3fff;
mem[890]<='h3fff;
mem[891]<='h3fff;
mem[892]<='h3fff;
mem[893]<='h3fff;
mem[894]<='h3fff;
mem[895]<='h3fff;
mem[896]<='h3fff;
mem[897]<='h3fff;
mem[898]<='h3fff;
mem[899]<='h3fff;
mem[900]<='h3fff;
mem[901]<='h3fff;
mem[902]<='h3fff;
mem[903]<='h3fff;
mem[904]<='h3fff;
mem[905]<='h3fff;
mem[906]<='h3fff;
mem[907]<='h3fff;
mem[908]<='h3fff;
mem[909]<='h3fff;
mem[910]<='h3fff;
mem[911]<='h3fff;
mem[912]<='h3fff;
mem[913]<='h1683;
mem[914]<='h0185;
mem[915]<='h0186;
mem[916]<='h2BB7;
mem[917]<='h3007;
mem[918]<='h1283;
mem[919]<='h0085;
mem[920]<='h30F9;
mem[921]<='h0086;
mem[922]<='h018C;
mem[923]<='h0A8C;
mem[924]<='h018D;
mem[925]<='h1283;
mem[926]<='h23B9;
mem[927]<='h300B;
mem[928]<='h0085;
mem[929]<='h0814;
mem[930]<='h0086;
mem[931]<='h018C;
mem[932]<='h0A8C;
mem[933]<='h018D;
mem[934]<='h23B9;
mem[935]<='h300D;
mem[936]<='h0085;
mem[937]<='h0815;
mem[938]<='h0086;
mem[939]<='h018C;
mem[940]<='h0A8C;
mem[941]<='h018D;
mem[942]<='h23B9;
mem[943]<='h300E;
mem[944]<='h0085;
mem[945]<='h0816;
mem[946]<='h0086;
mem[947]<='h018C;
mem[948]<='h0A8C;
mem[949]<='h018D;
mem[950]<='h23B9;
mem[951]<='h2B95;
mem[952]<='h2804;
mem[953]<='h080C;
mem[954]<='h008E;
mem[955]<='h080D;
mem[956]<='h008F;
mem[957]<='h080F;
mem[958]<='h040E;
mem[959]<='h1D03;
mem[960]<='h2BC2;
mem[961]<='h2BC3;
mem[962]<='h2BC4;
mem[963]<='h2BE5;
mem[964]<='h1283;
mem[965]<='h0190;
mem[966]<='h0A90;
mem[967]<='h0191;
mem[968]<='h0811;
mem[969]<='h0410;
mem[970]<='h1D03;
mem[971]<='h2BCD;
mem[972]<='h2BCE;
mem[973]<='h2BCF;
mem[974]<='h2BDA;
mem[975]<='h1283;
mem[976]<='h0890;
mem[977]<='h1903;
mem[978]<='h0391;
mem[979]<='h0390;
mem[980]<='h0811;
mem[981]<='h0410;
mem[982]<='h1D03;
mem[983]<='h2BD9;
mem[984]<='h2BDA;
mem[985]<='h2BCF;
mem[986]<='h1283;
mem[987]<='h088E;
mem[988]<='h1903;
mem[989]<='h038F;
mem[990]<='h038E;
mem[991]<='h080F;
mem[992]<='h040E;
mem[993]<='h1D03;
mem[994]<='h2BE4;
mem[995]<='h2BE5;
mem[996]<='h2BC4;
mem[997]<='h1283;
mem[998]<='h0008;
mem[999]<='h34C0;
mem[1000]<='h34F9;
mem[1001]<='h34A4;
mem[1002]<='h34B0;
mem[1003]<='h3499;
mem[1004]<='h3492;
mem[1005]<='h3482;
mem[1006]<='h34F8;
mem[1007]<='h3480;
mem[1008]<='h3490;
mem[1009]<='h3488;
mem[1010]<='h3483;
mem[1011]<='h34C6;
mem[1012]<='h34A1;
mem[1013]<='h3486;
mem[1014]<='h348E;
mem[1015]<='h3489;
mem[1016]<='h34C7;
mem[1017]<='h34C8;
mem[1018]<='h34C1;
mem[1019]<='h348C;
mem[1020]<='h34A3;
mem[1021]<='h34BF;
mem[1022]<='h34FF;
mem[1023]<='h34FF;








		end
	else
	begin
			if(en)
				OUT_DECODE<=mem[IN_PC];
			else
				OUT_DECODE<=OUT_DECODE;
	end
end
endmodule
		
