library verilog;
use verilog.vl_types.all;
entity memory is
    port(
        clock           : in     vl_logic;
        IN_PC           : in     vl_logic_vector(9 downto 0);
        en              : in     vl_logic;
        OUT_DECODE      : out    vl_logic_vector(13 downto 0)
    );
end memory;
